`default_nettype none

module tt_um_lif (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);
    // use bidirectionals as outputs
    //assign uio_oe = 8'b11111111;
    //assign uio_out[6:0] = 7'd0;
    //lif lif1(.current(ui_in), .clk(clk), .rst_n(rst_n), .spike(uio_out[7]), .state(uio_out));




    // lif lif2(.current(ui_in), .clk(clk), .rst_n(rst_n), .spike(uio_out[7]), .state(uio_out));

        // use bidirectionals as outputs
    assign uio_oe = 8'b11111111;

    // Default value for the 7 lower bits of uio_out
    assign uio_out[6:0] = 7'd0;

    wire spike;
    wire [7:0] state;
    wire [7:0] state_out;
    // Driving uo_out with state (example usage, modify as needed)
    assign uo_out = state;

    // Instantiate lif module
    lif lif1(
        .current(ui_in),
        .clk(clk),
        .rst_n(rst_n),
        .spike(spike),
        .state(state_out)
    );

    lif lif2(
        .current({uio_out[7], 7'b0000001}),
        .clk(clk),
        .rst_n(rst_n),
        .spike(uio_out[6]),
        .state(state)
    );

    // Assign spike to the highest bit of uio_out
    assign uio_out[7] = spike;

endmodule
